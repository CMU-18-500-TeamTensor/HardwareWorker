`ifndef MM_DEFINE
`define MM_DEFINE


typedef enum logic [5:0] {LINEAR, CONV, FLATTEN, MAXPOOL, RELU, SOFTMAX} layer_opcode;


`endif
