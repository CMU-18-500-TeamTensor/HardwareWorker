
module DPR();

endmodule: DPR

