`ifndef MM_DEFINE
`define MM_DEFINE

package MM_HANDSHAKE;

  parameter OPCODE_WIDTH;

endpackage: MM_HANDSHAKE

`endif
