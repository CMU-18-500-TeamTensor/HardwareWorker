
`ifndef TPP_OPCODE
`define TPP_OPCODE


typedef enum logic [31:0] {OP_ASN_MD=5, OP_ASN_DP=4, OP_M_FULL=6, OP_BATCH=8} tpp_opcode;

`endif
